/*
七段译码器

# 题目描述
七段显示译码器，可以把BCD码转换为七段显示码，从而可以显示数字0至数字9。
对应关系为：
0->0111111
1->0000110
2->1011011
3->1001111
4->1100110
5->1101101
6->1111101
7->0000111
8->1111111
9->1101111
其他输入->0000000
要求：在always块中使用if-else或case语句实现。

# 输入格式
输入为 din，为 4-bit wire。

# 输出格式
输出为 dout 从BCD转为七段显示码的结果，位宽为 7。
*/

module BCD7( 
    input [3:0] din, 
    output [6:0] dout
);
    reg [6:0] dout;
    always @(*)
    begin
        case(din)
            4'b0000: dout = 7'b0111111;
            4'b0001: dout = 7'b0000110;
            4'b0010: dout = 7'b1011011;
            4'b0011: dout = 7'b1001111;
            4'b0100: dout = 7'b1100110;
            4'b0101: dout = 7'b1101101;
            4'b0110: dout = 7'b1111101;
            4'b0111: dout = 7'b0000111;
            4'b1000: dout = 7'b1111111;
            4'b1001: dout = 7'b1101111;
            default: dout = 7'b0000000;
        endcase
    end
endmodule
