/*
输出1

# 题目描述
电路输出单比特信号1。

# 输入格式
无

# 输出格式
输出为out 位宽为1
*/

module One(
    output out
);
    assign out = 1'b1;
endmodule